`timescale 1ns / 1ps

module mul_top(input[3:0] x,y,
               input rst, go_mult, clk,
               output[7:0] product);

endmodule